/****************************************************************************
 * uex_sys_main.svh
 ****************************************************************************/

/**
 * Class: uex_sys_main
 * 
 * TODO: Add class documentation
 */
interface class uex_sys_main;

	pure virtual task main();

endclass


