/****************************************************************************
 * uex_sys_main.svh
 ****************************************************************************/

/**
 * Class: uex_sys_main
 * 
 * TODO: Add class documentation
 */
class uex_sys_main;

	virtual task main();
	endtask

endclass


