
`include "uvm_macros.svh"

package uex_ve_env_pkg;
	import uvm_pkg::*;
	import uex_pkg::*;

	`include "uex_ve_env.svh"
	
endpackage
