/****************************************************************************
 * uex_run_if.svh
 ****************************************************************************/

/**
 * Class: uex_run_if
 * 
 * TODO: Add class documentation
 */
interface class uex_run_if;

	pure virtual task run();

endclass


