/****************************************************************************
 * uex_c_thread.svh
 ****************************************************************************/

/**
 * Class: uex_c_thread
 * 
 * TODO: Add class documentation
 */
class uex_c_thread;

	function new();

	endfunction


endclass


