/****************************************************************************
 * uex_mem_services.svh
 ****************************************************************************/

/**
 * Class: uex_mem_services
 * 
 * TODO: Add class documentation
 */
interface class uex_mem_services extends uex_mem_access_services, uex_mem_alloc_services;

endclass


