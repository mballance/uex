/****************************************************************************
 * uex_ve_tb.sv
 ****************************************************************************/

/**
 * Module: uex_ve_tb
 * 
 * TODO: Add module documentation
 */
`include "uvm_macros.svh"
module uex_ve_tb;
	import uvm_pkg::*;
	import uex_ve_tests_pkg::*;
	
	initial begin
		run_test();
	end

endmodule

